`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer:        Tzu-Han Hsu
// Create Date:     07/29/2022 11:01:59 PM
// Module Name:     ZeroDetector_Group
// Project Name:    IEEE-754 & RISC-V Compatible Multiply-Accumulate Unit
// HDL(Version):    Verilog-2005
//
// Dependencies:    None
//
//////////////////////////////////////////////////////////////////////////////////
// Description:     Check if two groups are all zero
//
//////////////////////////////////////////////////////////////////////////////////
// Revision:
//
//////////////////////////////////////////////////////////////////////////////////


module ZeroDetector_Group #(
    parameter XLEN = 2
) (
    input [XLEN - 1 : 0] group_data_i,
    output group_zero_o );

    assign group_zero_o = &group_data_i;
    
endmodule